module arduino(in,lcdout);
input [3:0]in;
output [3:0]lcdout;
assign lcdout=in;
endmodule
